`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.02.2024 06:56:07
// Design Name: 
// Module Name: ieeeadd_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ieeeadd_tb( );
//wire [31:0] out;
//reg clk;
//reg [31:0] A,B;
//ieeedivision x1(out, A,B,clk);
//initial clk=1;
//always #10 clk=~clk;
//initial
//    begin
//     A=32'b0_10000011_00000000000000000000000;
//     B=32'b0_10000001_00000000000000000000000;
////    A=32'b0100_0000_0010_0000_0000_0000_0000_0000;
////    //B=32'b1011_1111_1100_0000_0000_0000_0000_0000;
////    B=0;
    
//   #20 
//   B=32'b0100_0000_0010_0000_0000_0000_0000_0000;
//   A=32'b0100_0000_0110_1100_1100_1100_1100_1101;
//    #20
////   //B=32'b0100_0000_0010_0000_0000_0000_0000_0000;
////   //B=32'b01000000101001100110011001100110; 
//   A=32'b0100_0000_0010_0000_0000_0000_0000_0000;
//    B=32'b1100_0001_0000_0100_1100_1100_1100_1101; 
//#20 
//A=32'b0_10000101_10010000000000000000000;
//B=32'b0_10000011_10010000000000000000000;
////    A = 32'b0_10000010_00111000000000000000000;
////        B = 32'b0_01111110_00100000000000000000000;
////  wire AEB,AGB,ALB;
////  reg clk;
////  reg [31:0]A,B;
////ieecomp x1(AEB,AGB,ALB,clk, A, B);
////initial clk=1;
////always #10 clk=~clk;
////initial
////    begin
////     A=32'b0_10000000_10000000000000000000000;
////     B=32'b0_10000000_10000000000000000000000;
//// #20
////    A=32'b1_10000000_00000000000000000000000;
////    B=32'b0_10000000_10000000000000000000000;
//// #20
////     A=32'b0_10000000_10000000000000000000000;
////     B=32'b0_10000000_10000000000000000000000;
//// #20
////     A=32'b0_10000000_00000000000000000000000;
////     B=32'b0_10000000_10000000000000000000000;
// #20
// A=32'b0_10000100_10010000000000000000000;
// B=32'b0_10000011_10010000000000000000000;
// #20
// A=32'b0_10000001_11100000000000000000000;
// B=32'b0_10000000_01000000000000000000000;
// #20
// A=32'b0_10000010_01000000000000000000000;
// B=32'b0_10000000_00000000000000000000000;
// #20
// A=32'b0_10000000_00000000000000000000000;
// B=32'b0_10000000_00000000000000000000000;
////     B=32'b0_10000000_00000000000000000000000;
////     A=32'b0_10000000_10000000000000000000000;
 reg clk;
 reg [31:0]A,B;
 reg [2:0] OPC;
wire [31:0] OUT;
wire  AEB,ALB,AGB;
FPU c1(clk, A,B,OPC,OUT,AEB, ALB,AGB);
initial clk=1;
always #20 clk=~clk;
initial
    begin
  OPC=5;
  A=32'b0_10000010_01001001100110011001101;
  B=32'b0_10000010_01001001100110011001101;
  #100
  OPC=0;
  A=32'b0_10000010_01001001100110011001101;
  B=32'b0_10000000_01011001100110011001101;
  #40
  OPC=1;
  A=32'b0_10000000_01000000000000000000000;
  B=32'b0_01111110_00000000000000000000000;
   #40
  OPC=2;
  A=32'b0_10000010_01000000000000000000000;
  B=32'b0_0111111000000000000000000000000;
  #40
  OPC=3;
  A=32'b0_10000000_11011001100110011001101;
  B=32'b0_10000000_01000000000000000000000;
  #40
  OPC=4;
 A=32'b0_10000000_01000000000000000000000;
 B=32'b0_10000000_01000000000000000000000;
 #40
 OPC=2;
  A=32'b0_10000010_01000000000000000000000;
  B=32'b0_0111111000000000000000000000000;
  
 #60 $finish;
    end
endmodule